module tfgrid