module vbuilder


