module base