module vbuilder
