module tfgrid
